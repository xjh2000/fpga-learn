module aes_sbox(input [7:0] in,    // input data byte
                output [7:0] out); // output data byte
    
    reg [7:0] Sbox[255:0];
    
    initial begin
        Sbox[0]   = 8'h63;
        Sbox[1]   = 8'h7c;
        Sbox[2]   = 8'h77;
        Sbox[3]   = 8'h7b;
        Sbox[4]   = 8'hf2;
        Sbox[5]   = 8'h6b;
        Sbox[6]   = 8'h6f;
        Sbox[7]   = 8'hc5;
        Sbox[8]   = 8'h30;
        Sbox[9]   = 8'h01;
        Sbox[10]  = 8'h67;
        Sbox[11]  = 8'h2b;
        Sbox[12]  = 8'hfe;
        Sbox[13]  = 8'hd7;
        Sbox[14]  = 8'hab;
        Sbox[15]  = 8'h76;
        Sbox[16]  = 8'hca;
        Sbox[17]  = 8'h82;
        Sbox[18]  = 8'hc9;
        Sbox[19]  = 8'h7d;
        Sbox[20]  = 8'hfa;
        Sbox[21]  = 8'h59;
        Sbox[22]  = 8'h47;
        Sbox[23]  = 8'hf0;
        Sbox[24]  = 8'had;
        Sbox[25]  = 8'hd4;
        Sbox[26]  = 8'ha2;
        Sbox[27]  = 8'haf;
        Sbox[28]  = 8'h9c;
        Sbox[29]  = 8'ha4;
        Sbox[30]  = 8'h72;
        Sbox[31]  = 8'hc0;
        Sbox[32]  = 8'hb7;
        Sbox[33]  = 8'hfd;
        Sbox[34]  = 8'h93;
        Sbox[35]  = 8'h26;
        Sbox[36]  = 8'h36;
        Sbox[37]  = 8'h3f;
        Sbox[38]  = 8'hf7;
        Sbox[39]  = 8'hcc;
        Sbox[40]  = 8'h34;
        Sbox[41]  = 8'ha5;
        Sbox[42]  = 8'he5;
        Sbox[43]  = 8'hf1;
        Sbox[44]  = 8'h71;
        Sbox[45]  = 8'hd8;
        Sbox[46]  = 8'h31;
        Sbox[47]  = 8'h15;
        Sbox[48]  = 8'h04;
        Sbox[49]  = 8'hc7;
        Sbox[50]  = 8'h23;
        Sbox[51]  = 8'hc3;
        Sbox[52]  = 8'h18;
        Sbox[53]  = 8'h96;
        Sbox[54]  = 8'h05;
        Sbox[55]  = 8'h9a;
        Sbox[56]  = 8'h07;
        Sbox[57]  = 8'h12;
        Sbox[58]  = 8'h80;
        Sbox[59]  = 8'he2;
        Sbox[60]  = 8'heb;
        Sbox[61]  = 8'h27;
        Sbox[62]  = 8'hb2;
        Sbox[63]  = 8'h75;
        Sbox[64]  = 8'h09;
        Sbox[65]  = 8'h83;
        Sbox[66]  = 8'h2c;
        Sbox[67]  = 8'h1a;
        Sbox[68]  = 8'h1b;
        Sbox[69]  = 8'h6e;
        Sbox[70]  = 8'h5a;
        Sbox[71]  = 8'ha0;
        Sbox[72]  = 8'h52;
        Sbox[73]  = 8'h3b;
        Sbox[74]  = 8'hd6;
        Sbox[75]  = 8'hb3;
        Sbox[76]  = 8'h29;
        Sbox[77]  = 8'he3;
        Sbox[78]  = 8'h2f;
        Sbox[79]  = 8'h84;
        Sbox[80]  = 8'h53;
        Sbox[81]  = 8'hd1;
        Sbox[82]  = 8'h00;
        Sbox[83]  = 8'hed;
        Sbox[84]  = 8'h20;
        Sbox[85]  = 8'hfc;
        Sbox[86]  = 8'hb1;
        Sbox[87]  = 8'h5b;
        Sbox[88]  = 8'h6a;
        Sbox[89]  = 8'hcb;
        Sbox[90]  = 8'hbe;
        Sbox[91]  = 8'h39;
        Sbox[92]  = 8'h4a;
        Sbox[93]  = 8'h4c;
        Sbox[94]  = 8'h58;
        Sbox[95]  = 8'hcf;
        Sbox[96]  = 8'hd0;
        Sbox[97]  = 8'hef;
        Sbox[98]  = 8'haa;
        Sbox[99]  = 8'hfb;
        Sbox[100] = 8'h43;
        Sbox[101] = 8'h4d;
        Sbox[102] = 8'h33;
        Sbox[103] = 8'h85;
        Sbox[104] = 8'h45;
        Sbox[105] = 8'hf9;
        Sbox[106] = 8'h02;
        Sbox[107] = 8'h7f;
        Sbox[108] = 8'h50;
        Sbox[109] = 8'h3c;
        Sbox[110] = 8'h9f;
        Sbox[111] = 8'ha8;
        Sbox[112] = 8'h51;
        Sbox[113] = 8'ha3;
        Sbox[114] = 8'h40;
        Sbox[115] = 8'h8f;
        Sbox[116] = 8'h92;
        Sbox[117] = 8'h9d;
        Sbox[118] = 8'h38;
        Sbox[119] = 8'hf5;
        Sbox[120] = 8'hbc;
        Sbox[121] = 8'hb6;
        Sbox[122] = 8'hda;
        Sbox[123] = 8'h21;
        Sbox[124] = 8'h10;
        Sbox[125] = 8'hff;
        Sbox[126] = 8'hf3;
        Sbox[127] = 8'hd2;
        Sbox[128] = 8'hcd;
        Sbox[129] = 8'h0c;
        Sbox[130] = 8'h13;
        Sbox[131] = 8'hec;
        Sbox[132] = 8'h5f;
        Sbox[133] = 8'h97;
        Sbox[134] = 8'h44;
        Sbox[135] = 8'h17;
        Sbox[136] = 8'hc4;
        Sbox[137] = 8'ha7;
        Sbox[138] = 8'h7e;
        Sbox[139] = 8'h3d;
        Sbox[140] = 8'h64;
        Sbox[141] = 8'h5d;
        Sbox[142] = 8'h19;
        Sbox[143] = 8'h73;
        Sbox[144] = 8'h60;
        Sbox[145] = 8'h81;
        Sbox[146] = 8'h4f;
        Sbox[147] = 8'hdc;
        Sbox[148] = 8'h22;
        Sbox[149] = 8'h2a;
        Sbox[150] = 8'h90;
        Sbox[151] = 8'h88;
        Sbox[152] = 8'h46;
        Sbox[153] = 8'hee;
        Sbox[154] = 8'hb8;
        Sbox[155] = 8'h14;
        Sbox[156] = 8'hde;
        Sbox[157] = 8'h5e;
        Sbox[158] = 8'h0b;
        Sbox[159] = 8'hdb;
        Sbox[160] = 8'he0;
        Sbox[161] = 8'h32;
        Sbox[162] = 8'h3a;
        Sbox[163] = 8'h0a;
        Sbox[164] = 8'h49;
        Sbox[165] = 8'h06;
        Sbox[166] = 8'h24;
        Sbox[167] = 8'h5c;
        Sbox[168] = 8'hc2;
        Sbox[169] = 8'hd3;
        Sbox[170] = 8'hac;
        Sbox[171] = 8'h62;
        Sbox[172] = 8'h91;
        Sbox[173] = 8'h95;
        Sbox[174] = 8'he4;
        Sbox[175] = 8'h79;
        Sbox[176] = 8'he7;
        Sbox[177] = 8'hc8;
        Sbox[178] = 8'h37;
        Sbox[179] = 8'h6d;
        Sbox[180] = 8'h8d;
        Sbox[181] = 8'hd5;
        Sbox[182] = 8'h4e;
        Sbox[183] = 8'ha9;
        Sbox[184] = 8'h6c;
        Sbox[185] = 8'h56;
        Sbox[186] = 8'hf4;
        Sbox[187] = 8'hea;
        Sbox[188] = 8'h65;
        Sbox[189] = 8'h7a;
        Sbox[190] = 8'hae;
        Sbox[191] = 8'h08;
        Sbox[192] = 8'hba;
        Sbox[193] = 8'h78;
        Sbox[194] = 8'h25;
        Sbox[195] = 8'h2e;
        Sbox[196] = 8'h1c;
        Sbox[197] = 8'ha6;
        Sbox[198] = 8'hb4;
        Sbox[199] = 8'hc6;
        Sbox[200] = 8'he8;
        Sbox[201] = 8'hdd;
        Sbox[202] = 8'h74;
        Sbox[203] = 8'h1f;
        Sbox[204] = 8'h4b;
        Sbox[205] = 8'hbd;
        Sbox[206] = 8'h8b;
        Sbox[207] = 8'h8a;
        Sbox[208] = 8'h70;
        Sbox[209] = 8'h3e;
        Sbox[210] = 8'hb5;
        Sbox[211] = 8'h66;
        Sbox[212] = 8'h48;
        Sbox[213] = 8'h03;
        Sbox[214] = 8'hf6;
        Sbox[215] = 8'h0e;
        Sbox[216] = 8'h61;
        Sbox[217] = 8'h35;
        Sbox[218] = 8'h57;
        Sbox[219] = 8'hb9;
        Sbox[220] = 8'h86;
        Sbox[221] = 8'hc1;
        Sbox[222] = 8'h1d;
        Sbox[223] = 8'h9e;
        Sbox[224] = 8'he1;
        Sbox[225] = 8'hf8;
        Sbox[226] = 8'h98;
        Sbox[227] = 8'h11;
        Sbox[228] = 8'h69;
        Sbox[229] = 8'hd9;
        Sbox[230] = 8'h8e;
        Sbox[231] = 8'h94;
        Sbox[232] = 8'h9b;
        Sbox[233] = 8'h1e;
        Sbox[234] = 8'h87;
        Sbox[235] = 8'he9;
        Sbox[236] = 8'hce;
        Sbox[237] = 8'h55;
        Sbox[238] = 8'h28;
        Sbox[239] = 8'hdf;
        Sbox[240] = 8'h8c;
        Sbox[241] = 8'ha1;
        Sbox[242] = 8'h89;
        Sbox[243] = 8'h0d;
        Sbox[244] = 8'hbf;
        Sbox[245] = 8'he6;
        Sbox[246] = 8'h42;
        Sbox[247] = 8'h68;
        Sbox[248] = 8'h41;
        Sbox[249] = 8'h99;
        Sbox[250] = 8'h2d;
        Sbox[251] = 8'h0f;
        Sbox[252] = 8'hb0;
        Sbox[253] = 8'h54;
        Sbox[254] = 8'hbb;
        Sbox[255] = 8'h16;
    end

    assign  out = Sbox[in];
    
endmodule
