//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:34:21 05/30/2021 
// Design Name: 
// Module Name:    fS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fS(W,rkey,w1);
  input[0:31] W;
  input[0:31] rkey;
  output[0:31] w1;
  wire[0:7] s[1:7];
 
 
  assign s[1]=~(W[16:23]);
  assign s[2]=(W[24:31]&s[1]);
  assign s[3]=(W[8:15]^W[0:7]);

  assign w1[16:23]=s[3]^s[2];
  assign s[4]=(W[0:7]|s[1]);
  assign s[5]=((W[24:31]^s[4]));

  assign w1[24:31]=W[8:15]^s[5];
  assign s[6]=(W[16:23]^W[8:15]);
  assign s[7]=(s[3]&s[6]);

  assign w1[8:15]=s[6]^s[7];
  assign w1[0:7]=((rkey[24:31]&rkey[16:23])&((~W[8:15]&~W[16:23])|(W[0:7]&~W[16:23]&~W[24:31])|(~W[0:7]&~W[16:23]&W[24:31])|(~W[0:7]&W[8:15]&W[16:23])))|
		 (((rkey[0:7]^rkey[8:15])&~rkey[24:31])&((~W[0:7]&~W[16:23]&W[24:31])|(~W[8:15]&W[16:23]&~W[24:31])|(W[0:7]&W[16:23]&W[24:31])|(W[0:7]&~W[8:15])))|
		 
		 ((~(rkey[0:7]^rkey[8:15])&~rkey[24:31])&((~W[8:15]&~W[24:31])|(~W[0:7]&~W[16:23]&~W[24:31])|(W[0:7]&~W[8:15]&~W[16:23])|(~W[0:7]&W[16:23]&W[24:31])))|
		
		 ((~rkey[16:23]&rkey[24:31])&((~W[0:7]&~W[16:23]&W[24:31])|(W[0:7]&W[16:23]&W[24:31])|(W[8:15]&W[16:23]&~W[24:31])|(W[0:7]&W[8:15])));
		 

 

endmodule